/ubc/ece/data/cmc2/kits/GPDK45/gsclib045_all_v4.4/gsclib045/lef/gsclib045_multibitsDFF.lef